module project(clk,rst_n,tx,in/*,in1,in2,in3,in4
,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14
,in15,in16*/,out/*,tt,l,o,oo*/);
input       clk/*,tt,l*/;
//input in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,in11,in12,in13,in14,in15,in16;

input       rst_n;
//output reg o,oo;
//reg[15:0] counter;

input [15:0] in;
output reg [15:0] out;
output      tx;
reg [7:0] code;
//reg write;
//reg w;
//u1 t(clk,0,code,tx);
/*always@(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,
in11,in12,in13,in14,in15,in16)
begin
if(in1)
begin
out<=16'b1111100110011111;
code<=8'b00000001;
end
else
if(in2)
begin
out<=16'b0010001000101111;
code<=8'b00000010;
end
else
if(in3)
begin
out<=16'b0000000000001111;
code<=8'b00000011;
end
else
if(in4)
begin
out<=16'b0001001001001000;
code<=8'b00000100;
end
else
if(in5)
begin
out<=16'b0100101010011000;
code<=8'b00000101;
end
else
if(in6)
begin
out<=16'b0000011001100000;
code<=8'b00000110;
end
else
if(in7)
begin
out<=16'b1110101011100000;
code<=8'b00000111;
end
else
if(in8)
begin
out<=16'b1000100010001000;
code<=8'b00001000;
end
else
if(in9)
begin
out<=16'b0000111110011111;
code<=8'b00001001;
end
else
if(in10)
begin
out<=16'b0101001001011000;
code<=8'b00001010;
end
else
if(in11)
begin
out<=16'b1001011001101001;
code<=8'b00001011;
end
else
if(in12)
begin
out<=16'b0000111100000000;
code<=8'b00001100;
end
else
if(in13)
begin
out<=16'b1111000100010001;
code<=8'b00001101;
end
else
if(in14)
begin
out<=16'b0010101001000010;
code<=8'b00001110;
end
else
if(in15)
begin
out<=16'b0100111111110100;
code<=8'b00001111;
end
else
if(in16)
begin
out<=16'b1000010000101111;
code<=8'b00010000;
end
else
begin
//out<=16'b0000000000000000;
//code<=8'b00000000;
end
end*/


/*always@(tt,l,w)
begin
if(w)
begin
write<=w;
end
if(~tt)
begin
o<=1'b0;
code=8'b00000011;
//write<=1;
end
else
begin
if(~l)
begin
oo<=1'b0;
code<=8'b00000010;
//write<=1;
end
else
begin
o<=1'b1;
oo<=1'b1;
code<=8'b00000000;
end
end
end*/


always@(in)
begin
case(in)

16'b0000000000000001:
begin //1
out<=16'b1111100110011111;
code<=8'b00000001; end
16'b0000000000000010:
begin//2
out<=16'b0010001000101111;
code<=8'b00000010;
end
16'b0000000000000100:
begin//3
out<=16'b0000000000001111;
code<=8'b00000011;
end
16'b0000000000001000:
begin//4
out<=16'b0000000000001111;
code<=8'b00000100;
end
16'b0000000000010000:
begin//5
out<=16'b0100101010011000;
code<=8'b00000101;
end
16'b0000000000100000:
begin//6
out<=16'b0000011001100000;
code<=8'b00000110;
end
16'b0000000001000000:
begin//7
out<=16'b1110101011100000;
code<=8'b00000111;
end
16'b0000000010000000:
begin//8
out<=16'b1000100010001000;
code<=8'b00001000;
end
16'b0000000100000000:
begin//9
out<=16'b0000111110011111;
code<=8'b00001001;
end
16'b0000001000000000:
begin//10
out<=16'b0101001001011000;
code<=8'b00001010;
end
16'b0000010000000000:
begin//11
out<=16'b1001011001101001;
code<=8'b00001011;
end
16'b0000100000000000:
begin//12
out<=16'b0000111100000000;
code<=8'b00001100;
end
16'b0001000000000000:
begin//13
out<=16'b1111000100010001;
code<=8'b00001101;
end
16'b0010000000000000:
begin//14
out<=16'b0010101001000010;
code<=8'b00001110;
end
16'b0100000000000000:
begin//15
out<=16'b0100111111110100;
code<=8'b00001111;
end
16'b1000000000000100:
begin
out<=16'b1000010000101111;
code<=8'b00010000;
end
default:begin
out<=16'b0000000000000000;
code<=8'b00000000;
end
endcase
end
/*always@(in1,in2,in3,in4,in5,in6,in7,in8,in9,in10,
in11,in12,in13,in14,in15,in16)
begin
if(in1)
begin
out<=16'b1111100110011111;
code<=8'b00000001;
end
else
begin
if(in2)
begin
out<=16'b0010001000101111;
code<=8'b00000010;
end
else
begin
if(in3)
begin
out<=16'b0000000000001111;
code<=8'b00000011;
end
else
begin
if(in4)
begin
out<=16'b0000000000001111;
code<=8'b00000011;
end
else
begin
if(in5)
begin
out<=16'b0100101010011000;
code<=8'b00000101;
end
else
begin
if(in6)
begin
out<=16'b0000011001100000;
code<=8'b00000110;
end
else
begin
if(in7)
begin
out<=16'b1110101011100000;
code<=8'b00000111;
end
else
begin
if(in8)
begin
out<=16'b1000100010001000;
code<=8'b00001000;
end
else
begin
if(in9)
begin
out<=16'b0000111110011111;
code<=8'b00001001;
end
else
begin
if(in10)
begin
out<=16'b0101001001011000;
code<=8'b00001010;
end
else
begin
if(in11)
begin
out<=16'b1001011001101001;
code<=8'b00001011;
end
else
begin
if(in12)
begin
out<=16'b0000111100000000;
code<=8'b00001100;
end
else
begin
if(in13)
begin
out<=16'b1111000100010001;
code<=8'b00001101;
end
else
begin
if(in14)
begin
out<=16'b0010101001000010;
code<=8'b00001110;
end
else
begin
if(in15)
begin
out<=16'b0100111111110100;
code<=8'b00001111;
end
else
begin
if(in16)
begin
out<=16'b1000010000101111;
code<=8'b00010000;
end
else
begin
out<=16'b0000000000000000;
//code<=8'b00000000;
end
end
end
end
end
end
end
end
end
end
end
end
end
end
end
end
end*/

u1 t(clk,0,code,tx);


endmodule
